module sine_lookup(index, out);
	input logic unsigned [9:0] index;
	output logic signed [23:0] out;
	always_comb begin
		case(index)
			0: out = 24'(0);
			1: out = 24'(51471);
			2: out = 24'(102941);
			3: out = 24'(154406);
			4: out = 24'(205866);
			5: out = 24'(257318);
			6: out = 24'(308761);
			7: out = 24'(360192);
			8: out = 24'(411609);
			9: out = 24'(463011);
			10: out = 24'(514395);
			11: out = 24'(565760);
			12: out = 24'(617104);
			13: out = 24'(668424);
			14: out = 24'(719720);
			15: out = 24'(770988);
			16: out = 24'(822227);
			17: out = 24'(873435);
			18: out = 24'(924610);
			19: out = 24'(975751);
			20: out = 24'(1026855);
			21: out = 24'(1077920);
			22: out = 24'(1128944);
			23: out = 24'(1179926);
			24: out = 24'(1230864);
			25: out = 24'(1281755);
			26: out = 24'(1332598);
			27: out = 24'(1383391);
			28: out = 24'(1434132);
			29: out = 24'(1484819);
			30: out = 24'(1535449);
			31: out = 24'(1586022);
			32: out = 24'(1636536);
			33: out = 24'(1686987);
			34: out = 24'(1737376);
			35: out = 24'(1787698);
			36: out = 24'(1837954);
			37: out = 24'(1888140);
			38: out = 24'(1938255);
			39: out = 24'(1988298);
			40: out = 24'(2038265);
			41: out = 24'(2088156);
			42: out = 24'(2137968);
			43: out = 24'(2187699);
			44: out = 24'(2237348);
			45: out = 24'(2286913);
			46: out = 24'(2336392);
			47: out = 24'(2385783);
			48: out = 24'(2435084);
			49: out = 24'(2484293);
			50: out = 24'(2533409);
			51: out = 24'(2582429);
			52: out = 24'(2631353);
			53: out = 24'(2680177);
			54: out = 24'(2728900);
			55: out = 24'(2777521);
			56: out = 24'(2826036);
			57: out = 24'(2874446);
			58: out = 24'(2922747);
			59: out = 24'(2970938);
			60: out = 24'(3019018);
			61: out = 24'(3066984);
			62: out = 24'(3114834);
			63: out = 24'(3162567);
			64: out = 24'(3210181);
			65: out = 24'(3257674);
			66: out = 24'(3305044);
			67: out = 24'(3352290);
			68: out = 24'(3399410);
			69: out = 24'(3446402);
			70: out = 24'(3493264);
			71: out = 24'(3539994);
			72: out = 24'(3586592);
			73: out = 24'(3633054);
			74: out = 24'(3679379);
			75: out = 24'(3725566);
			76: out = 24'(3771613);
			77: out = 24'(3817517);
			78: out = 24'(3863278);
			79: out = 24'(3908894);
			80: out = 24'(3954362);
			81: out = 24'(3999681);
			82: out = 24'(4044850);
			83: out = 24'(4089867);
			84: out = 24'(4134729);
			85: out = 24'(4179436);
			86: out = 24'(4223986);
			87: out = 24'(4268376);
			88: out = 24'(4312606);
			89: out = 24'(4356673);
			90: out = 24'(4400577);
			91: out = 24'(4444314);
			92: out = 24'(4487885);
			93: out = 24'(4531286);
			94: out = 24'(4574517);
			95: out = 24'(4617576);
			96: out = 24'(4660460);
			97: out = 24'(4703170);
			98: out = 24'(4745702);
			99: out = 24'(4788055);
			100: out = 24'(4830229);
			101: out = 24'(4872220);
			102: out = 24'(4914028);
			103: out = 24'(4955651);
			104: out = 24'(4997087);
			105: out = 24'(5038336);
			106: out = 24'(5079394);
			107: out = 24'(5120262);
			108: out = 24'(5160936);
			109: out = 24'(5201416);
			110: out = 24'(5241701);
			111: out = 24'(5281788);
			112: out = 24'(5321676);
			113: out = 24'(5361364);
			114: out = 24'(5400850);
			115: out = 24'(5440133);
			116: out = 24'(5479210);
			117: out = 24'(5518082);
			118: out = 24'(5556746);
			119: out = 24'(5595200);
			120: out = 24'(5633444);
			121: out = 24'(5671476);
			122: out = 24'(5709294);
			123: out = 24'(5746898);
			124: out = 24'(5784285);
			125: out = 24'(5821454);
			126: out = 24'(5858404);
			127: out = 24'(5895134);
			128: out = 24'(5931641);
			129: out = 24'(5967925);
			130: out = 24'(6003985);
			131: out = 24'(6039818);
			132: out = 24'(6075424);
			133: out = 24'(6110802);
			134: out = 24'(6145949);
			135: out = 24'(6180865);
			136: out = 24'(6215548);
			137: out = 24'(6249997);
			138: out = 24'(6284211);
			139: out = 24'(6318188);
			140: out = 24'(6351928);
			141: out = 24'(6385428);
			142: out = 24'(6418688);
			143: out = 24'(6451706);
			144: out = 24'(6484481);
			145: out = 24'(6517012);
			146: out = 24'(6549298);
			147: out = 24'(6581337);
			148: out = 24'(6613129);
			149: out = 24'(6644671);
			150: out = 24'(6675963);
			151: out = 24'(6707004);
			152: out = 24'(6737793);
			153: out = 24'(6768327);
			154: out = 24'(6798607);
			155: out = 24'(6828631);
			156: out = 24'(6858398);
			157: out = 24'(6887907);
			158: out = 24'(6917156);
			159: out = 24'(6946145);
			160: out = 24'(6974872);
			161: out = 24'(7003337);
			162: out = 24'(7031538);
			163: out = 24'(7059474);
			164: out = 24'(7087145);
			165: out = 24'(7114549);
			166: out = 24'(7141684);
			167: out = 24'(7168551);
			168: out = 24'(7195149);
			169: out = 24'(7221475);
			170: out = 24'(7247529);
			171: out = 24'(7273311);
			172: out = 24'(7298818);
			173: out = 24'(7324051);
			174: out = 24'(7349008);
			175: out = 24'(7373688);
			176: out = 24'(7398091);
			177: out = 24'(7422216);
			178: out = 24'(7446060);
			179: out = 24'(7469625);
			180: out = 24'(7492908);
			181: out = 24'(7515909);
			182: out = 24'(7538627);
			183: out = 24'(7561062);
			184: out = 24'(7583211);
			185: out = 24'(7605075);
			186: out = 24'(7626653);
			187: out = 24'(7647944);
			188: out = 24'(7668947);
			189: out = 24'(7689661);
			190: out = 24'(7710085);
			191: out = 24'(7730220);
			192: out = 24'(7750063);
			193: out = 24'(7769614);
			194: out = 24'(7788873);
			195: out = 24'(7807839);
			196: out = 24'(7826510);
			197: out = 24'(7844887);
			198: out = 24'(7862969);
			199: out = 24'(7880755);
			200: out = 24'(7898244);
			201: out = 24'(7915435);
			202: out = 24'(7932329);
			203: out = 24'(7948924);
			204: out = 24'(7965219);
			205: out = 24'(7981215);
			206: out = 24'(7996910);
			207: out = 24'(8012304);
			208: out = 24'(8027397);
			209: out = 24'(8042187);
			210: out = 24'(8056675);
			211: out = 24'(8070859);
			212: out = 24'(8084739);
			213: out = 24'(8098315);
			214: out = 24'(8111586);
			215: out = 24'(8124552);
			216: out = 24'(8137211);
			217: out = 24'(8149565);
			218: out = 24'(8161611);
			219: out = 24'(8173351);
			220: out = 24'(8184782);
			221: out = 24'(8195906);
			222: out = 24'(8206720);
			223: out = 24'(8217226);
			224: out = 24'(8227423);
			225: out = 24'(8237309);
			226: out = 24'(8246886);
			227: out = 24'(8256152);
			228: out = 24'(8265107);
			229: out = 24'(8273751);
			230: out = 24'(8282084);
			231: out = 24'(8290105);
			232: out = 24'(8297813);
			233: out = 24'(8305210);
			234: out = 24'(8312293);
			235: out = 24'(8319064);
			236: out = 24'(8325521);
			237: out = 24'(8331665);
			238: out = 24'(8337495);
			239: out = 24'(8343012);
			240: out = 24'(8348214);
			241: out = 24'(8353102);
			242: out = 24'(8357675);
			243: out = 24'(8361934);
			244: out = 24'(8365878);
			245: out = 24'(8369507);
			246: out = 24'(8372821);
			247: out = 24'(8375820);
			248: out = 24'(8378503);
			249: out = 24'(8380871);
			250: out = 24'(8382923);
			251: out = 24'(8384660);
			252: out = 24'(8386081);
			253: out = 24'(8387186);
			254: out = 24'(8387976);
			255: out = 24'(8388450);
			256: out = 24'(8388608);
			257: out = 24'(8388450);
			258: out = 24'(8387976);
			259: out = 24'(8387186);
			260: out = 24'(8386081);
			261: out = 24'(8384660);
			262: out = 24'(8382923);
			263: out = 24'(8380871);
			264: out = 24'(8378503);
			265: out = 24'(8375820);
			266: out = 24'(8372821);
			267: out = 24'(8369507);
			268: out = 24'(8365878);
			269: out = 24'(8361934);
			270: out = 24'(8357675);
			271: out = 24'(8353102);
			272: out = 24'(8348214);
			273: out = 24'(8343012);
			274: out = 24'(8337495);
			275: out = 24'(8331665);
			276: out = 24'(8325521);
			277: out = 24'(8319064);
			278: out = 24'(8312293);
			279: out = 24'(8305210);
			280: out = 24'(8297813);
			281: out = 24'(8290105);
			282: out = 24'(8282084);
			283: out = 24'(8273751);
			284: out = 24'(8265107);
			285: out = 24'(8256152);
			286: out = 24'(8246886);
			287: out = 24'(8237309);
			288: out = 24'(8227423);
			289: out = 24'(8217226);
			290: out = 24'(8206720);
			291: out = 24'(8195906);
			292: out = 24'(8184782);
			293: out = 24'(8173351);
			294: out = 24'(8161611);
			295: out = 24'(8149565);
			296: out = 24'(8137211);
			297: out = 24'(8124552);
			298: out = 24'(8111586);
			299: out = 24'(8098315);
			300: out = 24'(8084739);
			301: out = 24'(8070859);
			302: out = 24'(8056675);
			303: out = 24'(8042187);
			304: out = 24'(8027397);
			305: out = 24'(8012304);
			306: out = 24'(7996910);
			307: out = 24'(7981215);
			308: out = 24'(7965219);
			309: out = 24'(7948924);
			310: out = 24'(7932329);
			311: out = 24'(7915435);
			312: out = 24'(7898244);
			313: out = 24'(7880755);
			314: out = 24'(7862969);
			315: out = 24'(7844887);
			316: out = 24'(7826510);
			317: out = 24'(7807839);
			318: out = 24'(7788873);
			319: out = 24'(7769614);
			320: out = 24'(7750063);
			321: out = 24'(7730220);
			322: out = 24'(7710085);
			323: out = 24'(7689661);
			324: out = 24'(7668947);
			325: out = 24'(7647944);
			326: out = 24'(7626653);
			327: out = 24'(7605075);
			328: out = 24'(7583211);
			329: out = 24'(7561062);
			330: out = 24'(7538627);
			331: out = 24'(7515909);
			332: out = 24'(7492908);
			333: out = 24'(7469625);
			334: out = 24'(7446060);
			335: out = 24'(7422216);
			336: out = 24'(7398091);
			337: out = 24'(7373688);
			338: out = 24'(7349008);
			339: out = 24'(7324051);
			340: out = 24'(7298818);
			341: out = 24'(7273311);
			342: out = 24'(7247529);
			343: out = 24'(7221475);
			344: out = 24'(7195149);
			345: out = 24'(7168551);
			346: out = 24'(7141684);
			347: out = 24'(7114549);
			348: out = 24'(7087145);
			349: out = 24'(7059474);
			350: out = 24'(7031538);
			351: out = 24'(7003337);
			352: out = 24'(6974872);
			353: out = 24'(6946145);
			354: out = 24'(6917156);
			355: out = 24'(6887907);
			356: out = 24'(6858398);
			357: out = 24'(6828631);
			358: out = 24'(6798607);
			359: out = 24'(6768327);
			360: out = 24'(6737793);
			361: out = 24'(6707004);
			362: out = 24'(6675963);
			363: out = 24'(6644671);
			364: out = 24'(6613129);
			365: out = 24'(6581337);
			366: out = 24'(6549298);
			367: out = 24'(6517012);
			368: out = 24'(6484481);
			369: out = 24'(6451706);
			370: out = 24'(6418688);
			371: out = 24'(6385428);
			372: out = 24'(6351928);
			373: out = 24'(6318188);
			374: out = 24'(6284211);
			375: out = 24'(6249997);
			376: out = 24'(6215548);
			377: out = 24'(6180865);
			378: out = 24'(6145949);
			379: out = 24'(6110802);
			380: out = 24'(6075424);
			381: out = 24'(6039818);
			382: out = 24'(6003985);
			383: out = 24'(5967925);
			384: out = 24'(5931641);
			385: out = 24'(5895134);
			386: out = 24'(5858404);
			387: out = 24'(5821454);
			388: out = 24'(5784285);
			389: out = 24'(5746898);
			390: out = 24'(5709294);
			391: out = 24'(5671476);
			392: out = 24'(5633444);
			393: out = 24'(5595200);
			394: out = 24'(5556746);
			395: out = 24'(5518082);
			396: out = 24'(5479210);
			397: out = 24'(5440133);
			398: out = 24'(5400850);
			399: out = 24'(5361364);
			400: out = 24'(5321676);
			401: out = 24'(5281788);
			402: out = 24'(5241701);
			403: out = 24'(5201416);
			404: out = 24'(5160936);
			405: out = 24'(5120262);
			406: out = 24'(5079394);
			407: out = 24'(5038336);
			408: out = 24'(4997087);
			409: out = 24'(4955651);
			410: out = 24'(4914028);
			411: out = 24'(4872220);
			412: out = 24'(4830229);
			413: out = 24'(4788055);
			414: out = 24'(4745702);
			415: out = 24'(4703170);
			416: out = 24'(4660460);
			417: out = 24'(4617576);
			418: out = 24'(4574517);
			419: out = 24'(4531286);
			420: out = 24'(4487885);
			421: out = 24'(4444314);
			422: out = 24'(4400577);
			423: out = 24'(4356673);
			424: out = 24'(4312606);
			425: out = 24'(4268376);
			426: out = 24'(4223986);
			427: out = 24'(4179436);
			428: out = 24'(4134729);
			429: out = 24'(4089867);
			430: out = 24'(4044850);
			431: out = 24'(3999681);
			432: out = 24'(3954362);
			433: out = 24'(3908894);
			434: out = 24'(3863278);
			435: out = 24'(3817517);
			436: out = 24'(3771613);
			437: out = 24'(3725566);
			438: out = 24'(3679379);
			439: out = 24'(3633054);
			440: out = 24'(3586592);
			441: out = 24'(3539994);
			442: out = 24'(3493264);
			443: out = 24'(3446402);
			444: out = 24'(3399410);
			445: out = 24'(3352290);
			446: out = 24'(3305044);
			447: out = 24'(3257674);
			448: out = 24'(3210181);
			449: out = 24'(3162567);
			450: out = 24'(3114834);
			451: out = 24'(3066984);
			452: out = 24'(3019018);
			453: out = 24'(2970938);
			454: out = 24'(2922747);
			455: out = 24'(2874446);
			456: out = 24'(2826036);
			457: out = 24'(2777521);
			458: out = 24'(2728900);
			459: out = 24'(2680177);
			460: out = 24'(2631353);
			461: out = 24'(2582429);
			462: out = 24'(2533409);
			463: out = 24'(2484293);
			464: out = 24'(2435084);
			465: out = 24'(2385783);
			466: out = 24'(2336392);
			467: out = 24'(2286913);
			468: out = 24'(2237348);
			469: out = 24'(2187699);
			470: out = 24'(2137968);
			471: out = 24'(2088156);
			472: out = 24'(2038265);
			473: out = 24'(1988298);
			474: out = 24'(1938255);
			475: out = 24'(1888140);
			476: out = 24'(1837954);
			477: out = 24'(1787698);
			478: out = 24'(1737376);
			479: out = 24'(1686987);
			480: out = 24'(1636536);
			481: out = 24'(1586022);
			482: out = 24'(1535449);
			483: out = 24'(1484819);
			484: out = 24'(1434132);
			485: out = 24'(1383391);
			486: out = 24'(1332598);
			487: out = 24'(1281755);
			488: out = 24'(1230864);
			489: out = 24'(1179926);
			490: out = 24'(1128944);
			491: out = 24'(1077920);
			492: out = 24'(1026855);
			493: out = 24'(975751);
			494: out = 24'(924610);
			495: out = 24'(873435);
			496: out = 24'(822227);
			497: out = 24'(770988);
			498: out = 24'(719720);
			499: out = 24'(668424);
			500: out = 24'(617104);
			501: out = 24'(565760);
			502: out = 24'(514395);
			503: out = 24'(463011);
			504: out = 24'(411609);
			505: out = 24'(360192);
			506: out = 24'(308761);
			507: out = 24'(257318);
			508: out = 24'(205866);
			509: out = 24'(154406);
			510: out = 24'(102941);
			511: out = 24'(51471);
			512: out = 24'(0);
			513: out = 24'(-51471);
			514: out = 24'(-102941);
			515: out = 24'(-154406);
			516: out = 24'(-205866);
			517: out = 24'(-257318);
			518: out = 24'(-308761);
			519: out = 24'(-360192);
			520: out = 24'(-411609);
			521: out = 24'(-463011);
			522: out = 24'(-514395);
			523: out = 24'(-565760);
			524: out = 24'(-617104);
			525: out = 24'(-668424);
			526: out = 24'(-719720);
			527: out = 24'(-770988);
			528: out = 24'(-822227);
			529: out = 24'(-873435);
			530: out = 24'(-924610);
			531: out = 24'(-975751);
			532: out = 24'(-1026855);
			533: out = 24'(-1077920);
			534: out = 24'(-1128944);
			535: out = 24'(-1179926);
			536: out = 24'(-1230864);
			537: out = 24'(-1281755);
			538: out = 24'(-1332598);
			539: out = 24'(-1383391);
			540: out = 24'(-1434132);
			541: out = 24'(-1484819);
			542: out = 24'(-1535449);
			543: out = 24'(-1586022);
			544: out = 24'(-1636536);
			545: out = 24'(-1686987);
			546: out = 24'(-1737376);
			547: out = 24'(-1787698);
			548: out = 24'(-1837954);
			549: out = 24'(-1888140);
			550: out = 24'(-1938255);
			551: out = 24'(-1988298);
			552: out = 24'(-2038265);
			553: out = 24'(-2088156);
			554: out = 24'(-2137968);
			555: out = 24'(-2187699);
			556: out = 24'(-2237348);
			557: out = 24'(-2286913);
			558: out = 24'(-2336392);
			559: out = 24'(-2385783);
			560: out = 24'(-2435084);
			561: out = 24'(-2484293);
			562: out = 24'(-2533409);
			563: out = 24'(-2582429);
			564: out = 24'(-2631353);
			565: out = 24'(-2680177);
			566: out = 24'(-2728900);
			567: out = 24'(-2777521);
			568: out = 24'(-2826036);
			569: out = 24'(-2874446);
			570: out = 24'(-2922747);
			571: out = 24'(-2970938);
			572: out = 24'(-3019018);
			573: out = 24'(-3066984);
			574: out = 24'(-3114834);
			575: out = 24'(-3162567);
			576: out = 24'(-3210181);
			577: out = 24'(-3257674);
			578: out = 24'(-3305044);
			579: out = 24'(-3352290);
			580: out = 24'(-3399410);
			581: out = 24'(-3446402);
			582: out = 24'(-3493264);
			583: out = 24'(-3539994);
			584: out = 24'(-3586592);
			585: out = 24'(-3633054);
			586: out = 24'(-3679379);
			587: out = 24'(-3725566);
			588: out = 24'(-3771613);
			589: out = 24'(-3817517);
			590: out = 24'(-3863278);
			591: out = 24'(-3908894);
			592: out = 24'(-3954362);
			593: out = 24'(-3999681);
			594: out = 24'(-4044850);
			595: out = 24'(-4089867);
			596: out = 24'(-4134729);
			597: out = 24'(-4179436);
			598: out = 24'(-4223986);
			599: out = 24'(-4268376);
			600: out = 24'(-4312606);
			601: out = 24'(-4356673);
			602: out = 24'(-4400577);
			603: out = 24'(-4444314);
			604: out = 24'(-4487885);
			605: out = 24'(-4531286);
			606: out = 24'(-4574517);
			607: out = 24'(-4617576);
			608: out = 24'(-4660460);
			609: out = 24'(-4703170);
			610: out = 24'(-4745702);
			611: out = 24'(-4788055);
			612: out = 24'(-4830229);
			613: out = 24'(-4872220);
			614: out = 24'(-4914028);
			615: out = 24'(-4955651);
			616: out = 24'(-4997087);
			617: out = 24'(-5038336);
			618: out = 24'(-5079394);
			619: out = 24'(-5120262);
			620: out = 24'(-5160936);
			621: out = 24'(-5201416);
			622: out = 24'(-5241701);
			623: out = 24'(-5281788);
			624: out = 24'(-5321676);
			625: out = 24'(-5361364);
			626: out = 24'(-5400850);
			627: out = 24'(-5440133);
			628: out = 24'(-5479210);
			629: out = 24'(-5518082);
			630: out = 24'(-5556746);
			631: out = 24'(-5595200);
			632: out = 24'(-5633444);
			633: out = 24'(-5671476);
			634: out = 24'(-5709294);
			635: out = 24'(-5746898);
			636: out = 24'(-5784285);
			637: out = 24'(-5821454);
			638: out = 24'(-5858404);
			639: out = 24'(-5895134);
			640: out = 24'(-5931641);
			641: out = 24'(-5967925);
			642: out = 24'(-6003985);
			643: out = 24'(-6039818);
			644: out = 24'(-6075424);
			645: out = 24'(-6110802);
			646: out = 24'(-6145949);
			647: out = 24'(-6180865);
			648: out = 24'(-6215548);
			649: out = 24'(-6249997);
			650: out = 24'(-6284211);
			651: out = 24'(-6318188);
			652: out = 24'(-6351928);
			653: out = 24'(-6385428);
			654: out = 24'(-6418688);
			655: out = 24'(-6451706);
			656: out = 24'(-6484481);
			657: out = 24'(-6517012);
			658: out = 24'(-6549298);
			659: out = 24'(-6581337);
			660: out = 24'(-6613129);
			661: out = 24'(-6644671);
			662: out = 24'(-6675963);
			663: out = 24'(-6707004);
			664: out = 24'(-6737793);
			665: out = 24'(-6768327);
			666: out = 24'(-6798607);
			667: out = 24'(-6828631);
			668: out = 24'(-6858398);
			669: out = 24'(-6887907);
			670: out = 24'(-6917156);
			671: out = 24'(-6946145);
			672: out = 24'(-6974872);
			673: out = 24'(-7003337);
			674: out = 24'(-7031538);
			675: out = 24'(-7059474);
			676: out = 24'(-7087145);
			677: out = 24'(-7114549);
			678: out = 24'(-7141684);
			679: out = 24'(-7168551);
			680: out = 24'(-7195149);
			681: out = 24'(-7221475);
			682: out = 24'(-7247529);
			683: out = 24'(-7273311);
			684: out = 24'(-7298818);
			685: out = 24'(-7324051);
			686: out = 24'(-7349008);
			687: out = 24'(-7373688);
			688: out = 24'(-7398091);
			689: out = 24'(-7422216);
			690: out = 24'(-7446060);
			691: out = 24'(-7469625);
			692: out = 24'(-7492908);
			693: out = 24'(-7515909);
			694: out = 24'(-7538627);
			695: out = 24'(-7561062);
			696: out = 24'(-7583211);
			697: out = 24'(-7605075);
			698: out = 24'(-7626653);
			699: out = 24'(-7647944);
			700: out = 24'(-7668947);
			701: out = 24'(-7689661);
			702: out = 24'(-7710085);
			703: out = 24'(-7730220);
			704: out = 24'(-7750063);
			705: out = 24'(-7769614);
			706: out = 24'(-7788873);
			707: out = 24'(-7807839);
			708: out = 24'(-7826510);
			709: out = 24'(-7844887);
			710: out = 24'(-7862969);
			711: out = 24'(-7880755);
			712: out = 24'(-7898244);
			713: out = 24'(-7915435);
			714: out = 24'(-7932329);
			715: out = 24'(-7948924);
			716: out = 24'(-7965219);
			717: out = 24'(-7981215);
			718: out = 24'(-7996910);
			719: out = 24'(-8012304);
			720: out = 24'(-8027397);
			721: out = 24'(-8042187);
			722: out = 24'(-8056675);
			723: out = 24'(-8070859);
			724: out = 24'(-8084739);
			725: out = 24'(-8098315);
			726: out = 24'(-8111586);
			727: out = 24'(-8124552);
			728: out = 24'(-8137211);
			729: out = 24'(-8149565);
			730: out = 24'(-8161611);
			731: out = 24'(-8173351);
			732: out = 24'(-8184782);
			733: out = 24'(-8195906);
			734: out = 24'(-8206720);
			735: out = 24'(-8217226);
			736: out = 24'(-8227423);
			737: out = 24'(-8237309);
			738: out = 24'(-8246886);
			739: out = 24'(-8256152);
			740: out = 24'(-8265107);
			741: out = 24'(-8273751);
			742: out = 24'(-8282084);
			743: out = 24'(-8290105);
			744: out = 24'(-8297813);
			745: out = 24'(-8305210);
			746: out = 24'(-8312293);
			747: out = 24'(-8319064);
			748: out = 24'(-8325521);
			749: out = 24'(-8331665);
			750: out = 24'(-8337495);
			751: out = 24'(-8343012);
			752: out = 24'(-8348214);
			753: out = 24'(-8353102);
			754: out = 24'(-8357675);
			755: out = 24'(-8361934);
			756: out = 24'(-8365878);
			757: out = 24'(-8369507);
			758: out = 24'(-8372821);
			759: out = 24'(-8375820);
			760: out = 24'(-8378503);
			761: out = 24'(-8380871);
			762: out = 24'(-8382923);
			763: out = 24'(-8384660);
			764: out = 24'(-8386081);
			765: out = 24'(-8387186);
			766: out = 24'(-8387976);
			767: out = 24'(-8388450);
			768: out = 24'(-8388608);
			769: out = 24'(-8388450);
			770: out = 24'(-8387976);
			771: out = 24'(-8387186);
			772: out = 24'(-8386081);
			773: out = 24'(-8384660);
			774: out = 24'(-8382923);
			775: out = 24'(-8380871);
			776: out = 24'(-8378503);
			777: out = 24'(-8375820);
			778: out = 24'(-8372821);
			779: out = 24'(-8369507);
			780: out = 24'(-8365878);
			781: out = 24'(-8361934);
			782: out = 24'(-8357675);
			783: out = 24'(-8353102);
			784: out = 24'(-8348214);
			785: out = 24'(-8343012);
			786: out = 24'(-8337495);
			787: out = 24'(-8331665);
			788: out = 24'(-8325521);
			789: out = 24'(-8319064);
			790: out = 24'(-8312293);
			791: out = 24'(-8305210);
			792: out = 24'(-8297813);
			793: out = 24'(-8290105);
			794: out = 24'(-8282084);
			795: out = 24'(-8273751);
			796: out = 24'(-8265107);
			797: out = 24'(-8256152);
			798: out = 24'(-8246886);
			799: out = 24'(-8237309);
			800: out = 24'(-8227423);
			801: out = 24'(-8217226);
			802: out = 24'(-8206720);
			803: out = 24'(-8195906);
			804: out = 24'(-8184782);
			805: out = 24'(-8173351);
			806: out = 24'(-8161611);
			807: out = 24'(-8149565);
			808: out = 24'(-8137211);
			809: out = 24'(-8124552);
			810: out = 24'(-8111586);
			811: out = 24'(-8098315);
			812: out = 24'(-8084739);
			813: out = 24'(-8070859);
			814: out = 24'(-8056675);
			815: out = 24'(-8042187);
			816: out = 24'(-8027397);
			817: out = 24'(-8012304);
			818: out = 24'(-7996910);
			819: out = 24'(-7981215);
			820: out = 24'(-7965219);
			821: out = 24'(-7948924);
			822: out = 24'(-7932329);
			823: out = 24'(-7915435);
			824: out = 24'(-7898244);
			825: out = 24'(-7880755);
			826: out = 24'(-7862969);
			827: out = 24'(-7844887);
			828: out = 24'(-7826510);
			829: out = 24'(-7807839);
			830: out = 24'(-7788873);
			831: out = 24'(-7769614);
			832: out = 24'(-7750063);
			833: out = 24'(-7730220);
			834: out = 24'(-7710085);
			835: out = 24'(-7689661);
			836: out = 24'(-7668947);
			837: out = 24'(-7647944);
			838: out = 24'(-7626653);
			839: out = 24'(-7605075);
			840: out = 24'(-7583211);
			841: out = 24'(-7561062);
			842: out = 24'(-7538627);
			843: out = 24'(-7515909);
			844: out = 24'(-7492908);
			845: out = 24'(-7469625);
			846: out = 24'(-7446060);
			847: out = 24'(-7422216);
			848: out = 24'(-7398091);
			849: out = 24'(-7373688);
			850: out = 24'(-7349008);
			851: out = 24'(-7324051);
			852: out = 24'(-7298818);
			853: out = 24'(-7273311);
			854: out = 24'(-7247529);
			855: out = 24'(-7221475);
			856: out = 24'(-7195149);
			857: out = 24'(-7168551);
			858: out = 24'(-7141684);
			859: out = 24'(-7114549);
			860: out = 24'(-7087145);
			861: out = 24'(-7059474);
			862: out = 24'(-7031538);
			863: out = 24'(-7003337);
			864: out = 24'(-6974872);
			865: out = 24'(-6946145);
			866: out = 24'(-6917156);
			867: out = 24'(-6887907);
			868: out = 24'(-6858398);
			869: out = 24'(-6828631);
			870: out = 24'(-6798607);
			871: out = 24'(-6768327);
			872: out = 24'(-6737793);
			873: out = 24'(-6707004);
			874: out = 24'(-6675963);
			875: out = 24'(-6644671);
			876: out = 24'(-6613129);
			877: out = 24'(-6581337);
			878: out = 24'(-6549298);
			879: out = 24'(-6517012);
			880: out = 24'(-6484481);
			881: out = 24'(-6451706);
			882: out = 24'(-6418688);
			883: out = 24'(-6385428);
			884: out = 24'(-6351928);
			885: out = 24'(-6318188);
			886: out = 24'(-6284211);
			887: out = 24'(-6249997);
			888: out = 24'(-6215548);
			889: out = 24'(-6180865);
			890: out = 24'(-6145949);
			891: out = 24'(-6110802);
			892: out = 24'(-6075424);
			893: out = 24'(-6039818);
			894: out = 24'(-6003985);
			895: out = 24'(-5967925);
			896: out = 24'(-5931641);
			897: out = 24'(-5895134);
			898: out = 24'(-5858404);
			899: out = 24'(-5821454);
			900: out = 24'(-5784285);
			901: out = 24'(-5746898);
			902: out = 24'(-5709294);
			903: out = 24'(-5671476);
			904: out = 24'(-5633444);
			905: out = 24'(-5595200);
			906: out = 24'(-5556746);
			907: out = 24'(-5518082);
			908: out = 24'(-5479210);
			909: out = 24'(-5440133);
			910: out = 24'(-5400850);
			911: out = 24'(-5361364);
			912: out = 24'(-5321676);
			913: out = 24'(-5281788);
			914: out = 24'(-5241701);
			915: out = 24'(-5201416);
			916: out = 24'(-5160936);
			917: out = 24'(-5120262);
			918: out = 24'(-5079394);
			919: out = 24'(-5038336);
			920: out = 24'(-4997087);
			921: out = 24'(-4955651);
			922: out = 24'(-4914028);
			923: out = 24'(-4872220);
			924: out = 24'(-4830229);
			925: out = 24'(-4788055);
			926: out = 24'(-4745702);
			927: out = 24'(-4703170);
			928: out = 24'(-4660460);
			929: out = 24'(-4617576);
			930: out = 24'(-4574517);
			931: out = 24'(-4531286);
			932: out = 24'(-4487885);
			933: out = 24'(-4444314);
			934: out = 24'(-4400577);
			935: out = 24'(-4356673);
			936: out = 24'(-4312606);
			937: out = 24'(-4268376);
			938: out = 24'(-4223986);
			939: out = 24'(-4179436);
			940: out = 24'(-4134729);
			941: out = 24'(-4089867);
			942: out = 24'(-4044850);
			943: out = 24'(-3999681);
			944: out = 24'(-3954362);
			945: out = 24'(-3908894);
			946: out = 24'(-3863278);
			947: out = 24'(-3817517);
			948: out = 24'(-3771613);
			949: out = 24'(-3725566);
			950: out = 24'(-3679379);
			951: out = 24'(-3633054);
			952: out = 24'(-3586592);
			953: out = 24'(-3539994);
			954: out = 24'(-3493264);
			955: out = 24'(-3446402);
			956: out = 24'(-3399410);
			957: out = 24'(-3352290);
			958: out = 24'(-3305044);
			959: out = 24'(-3257674);
			960: out = 24'(-3210181);
			961: out = 24'(-3162567);
			962: out = 24'(-3114834);
			963: out = 24'(-3066984);
			964: out = 24'(-3019018);
			965: out = 24'(-2970938);
			966: out = 24'(-2922747);
			967: out = 24'(-2874446);
			968: out = 24'(-2826036);
			969: out = 24'(-2777521);
			970: out = 24'(-2728900);
			971: out = 24'(-2680177);
			972: out = 24'(-2631353);
			973: out = 24'(-2582429);
			974: out = 24'(-2533409);
			975: out = 24'(-2484293);
			976: out = 24'(-2435084);
			977: out = 24'(-2385783);
			978: out = 24'(-2336392);
			979: out = 24'(-2286913);
			980: out = 24'(-2237348);
			981: out = 24'(-2187699);
			982: out = 24'(-2137968);
			983: out = 24'(-2088156);
			984: out = 24'(-2038265);
			985: out = 24'(-1988298);
			986: out = 24'(-1938255);
			987: out = 24'(-1888140);
			988: out = 24'(-1837954);
			989: out = 24'(-1787698);
			990: out = 24'(-1737376);
			991: out = 24'(-1686987);
			992: out = 24'(-1636536);
			993: out = 24'(-1586022);
			994: out = 24'(-1535449);
			995: out = 24'(-1484819);
			996: out = 24'(-1434132);
			997: out = 24'(-1383391);
			998: out = 24'(-1332598);
			999: out = 24'(-1281755);
			1000: out = 24'(-1230864);
			1001: out = 24'(-1179926);
			1002: out = 24'(-1128944);
			1003: out = 24'(-1077920);
			1004: out = 24'(-1026855);
			1005: out = 24'(-975751);
			1006: out = 24'(-924610);
			1007: out = 24'(-873435);
			1008: out = 24'(-822227);
			1009: out = 24'(-770988);
			1010: out = 24'(-719720);
			1011: out = 24'(-668424);
			1012: out = 24'(-617104);
			1013: out = 24'(-565760);
			1014: out = 24'(-514395);
			1015: out = 24'(-463011);
			1016: out = 24'(-411609);
			1017: out = 24'(-360192);
			1018: out = 24'(-308761);
			1019: out = 24'(-257318);
			1020: out = 24'(-205866);
			1021: out = 24'(-154406);
			1022: out = 24'(-102941);
			1023: out = 24'(-51471);
			default: out = 24'(0);
		endcase
	end
endmodule
